
module fp_multiplier_tb;

reg[31:0] a;
reg[31:0] b;
wire[31:0] result;

fp_multiplier FPA(.a(a), .b(b), .result(result));

initial begin
	a <= 32'b10111111100010000000000000000000;
	b <= 32'b11000000011001000000000000000000;
	#60
	a <= 32'b01000001001101000001111010111000;
	b <= 32'b11000001010101000000000000000000;
	#60
	a <= 32'b01000001110001100000000000000000;
	b <= 32'b01000001110001100000000000000000;
	#60
	a <= 32'b11000010101110010000000000000000;
	b <= 32'b01000010100111011000000000000000;
end

endmodule