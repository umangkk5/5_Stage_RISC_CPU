
module fp_adder_tb;

reg[31:0] a;
reg[31:0] b;
wire[31:0] result;

fp_adder FPA(.a(a), .b(b), .result(result));

initial begin
	a <= 32'b01000001100000000000000000001100;
	b <= 32'b01010001100011000000000000000000;
	#60
	a <= 32'b01000000010100000000000000000000;
	b <= 32'b00111111110000000000000000000000;
	#60
	a <= 32'b11000001110001000000000000000000;
	b <= 32'b01000001110011100000000000000000;
	#60
	a <= 32'b11000001110001000000000000000000;
	b <= 32'b11000001110011100000000000000000;
end

endmodule